library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity ioport is
	 Generic (BASE_ADDR	: integer := 16#19#);
    Port ( clk : in  STD_LOGIC;
	       Rst : in  STD_LOGIC;
           addr : in  STD_LOGIC_VECTOR (5 downto 0);
           ioread : out  STD_LOGIC_VECTOR (7 downto 0);
           iowrite : in  STD_LOGIC_VECTOR (7 downto 0);
           rd : in  STD_LOGIC;
           wr : in  STD_LOGIC;
		   ioport : inout  STD_LOGIC_VECTOR (7 downto 0));
end ioport;

architecture ioport_architecture of ioport is

constant PORT_ADDR : integer := BASE_ADDR + 2;
constant DDR_ADDR : integer := BASE_ADDR + 1;
constant PIN_ADDR : integer := BASE_ADDR;

signal port_reg, pin_reg, ddr_reg: std_logic_vector(7 downto 0);


begin

  proc : process(clk,Rst)
    variable adr_int : natural;
    -- variable rdwr : std_logic_vector(1 downto 0);

  begin

    if Rst = '1' then
      port_reg <= (others =>'Z');
      ddr_reg <= (others =>'0');
      pin_reg <= (others => '0');

    elsif rising_edge(clk) then
      adr_int := CONV_INTEGER(unsigned(addr));
      -- rdwr := rd & wr;

      if addr = PORT_ADDR then
            port_reg <= iowrite;
      elsif addr = DDR_ADDR then
            ddr_reg <= iowrite;
      elsif addr = PIN_ADDR then
            ioread <= pin_reg;
      end if;

      bits_port : for i in 0 to 7 loop
        if ddr_reg(i) = '0' then
          port_reg(i) <= 'Z';
        end if;
      end loop;

      read_write : for i in 0 to 7 loop
        if ddr_reg(i) = '1' then --sortie
          ioport(i) <= port_reg(i);
          pin_reg(i) <= '0';
        elsif ddr_reg(i) = '0' then --entrée
          pin_reg(i) <= ioport(i);
        end if;
      end loop;
    end if;
  end process;

end ioport_architecture;

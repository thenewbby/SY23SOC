-- filename : build/pm.hex
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity pm is
	Port (
           clk    : in std_logic;
           PM_A   : in std_logic_vector(15 downto 0);
           PM_Drd : out std_logic_vector(15 downto 0));
end pm;

architecture Arch of pm is

-- datas
type PM_mem_type is array(0 to 4095) of std_logic_vector(15 downto 0);
signal PM_mem : PM_mem_type := (
    x"C012", x"C019", x"C018", x"C017", x"C016", x"C015", x"C014", x"C013", 
    x"C012", x"C011", x"C010", x"C00F", x"C00E", x"C00D", x"C00C", x"C00B", 
    x"C00A", x"C009", x"C008", x"2411", x"BE1F", x"E5CF", x"E0D2", x"BFDE", 
    x"BFCD", x"D002", x"C008", x"CFE4", x"E880", x"BD8D", x"E182", x"BD8F", 
    x"E482", x"BF80", x"CFFF", x"94F8", x"CFFF", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", 
    x"0000", x"0000", x"0000" );
-- program size 74 / 4096

begin

   pmproc : process (clk)
     variable a_int : natural;
   begin
     if (clk'event and clk='1') then
        a_int := CONV_INTEGER(PM_A);
        PM_Drd <= PM_mem(a_int);
     end if;
  end process pmproc;

end architecture Arch;

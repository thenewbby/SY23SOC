--test bench file for prediviseur component
